module simplest(input i, output o);
    assign o = i;
endmodule